// Muhammad Tahir Zia 
// 2021465

`timescale 1ns/1ps

module multiply6bits_tb;
reg [5:0] inp1, inp2;
wire [11:0] product;
  
multiply6bits uut (.product(product),.inp1(inp1),.inp2(inp2));
  
initial begin
inp1 = 0; inp2 = 0;
#10;
    
inp1 = 6'b101010; inp2 = 6'b101000;
#10;
    
inp1 = 6'b101011; inp2 = 6'b101010;
#10;
    
inp1 = 6'b101011; inp2 = 6'b101100;
#10;
    
inp1 = 6'b101000; inp2 = 6'b100000;
#10;
    
$finish;
end
  
initial begin
$monitor("Time=%0t inp1=%d inp2=%d product=%d expected=%d", 
$time, inp1, inp2, product, inp1*inp2);
end
  
endmodule